architecture archRTL of cy_mxs40_tcpwm_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_dw_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_gpio_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_smartio_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_smif_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_ble_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_scb_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_scb_v1_10 is
begin
end archRTL;

architecture archRTL of cy_mxs40_csd_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_usb_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_ipc_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_crypto_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_profile_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_i2s_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_pdm_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_lpcomp_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_isr_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_samplehold_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_csidac_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_opamp_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_lcd_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_ctdac_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_ctdac_v1_10 is
begin
end archRTL;

architecture archRTL of cy_mxs40_sar_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_sarmux_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_temp_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_mcwdt_v1_0 is
begin
end archRTL;

architecture archRTL of cy_mxs40_rtc_v1_0 is
begin
end archRTL;
