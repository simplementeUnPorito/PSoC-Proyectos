-- cy_psoc3.vhp
--

--------------------------------------------------------------------------------
-- PSoC3 Component Declarations
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
package psoc3pkg is

-- PSoC3 Components
component cy_psoc3_dp8
    generic(cy_dpconfig_a : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     ce0_sync : std_logic := '1';
     cl0_sync : std_logic := '1';
     z0_sync : std_logic := '1';
     ff0_sync : std_logic := '1';
     ce1_sync : std_logic := '1';
     cl1_sync : std_logic := '1';
     z1_sync : std_logic := '1';
     ff1_sync : std_logic := '1';
     ov_msb_sync : std_logic := '1';
     co_msb_sync : std_logic := '1';
     cmsb_sync : std_logic := '1';
     so_sync : std_logic := '1';
     f0_bus_sync : std_logic := '1';
     f0_blk_sync : std_logic := '1';
     f1_bus_sync : std_logic := '1';
     f1_blk_sync : std_logic := '1');
    port ( reset : in std_logic := '0';
     clk : in std_logic;
     cs_addr : in std_logic_vector (2 downto 0);
     route_si : in std_logic;
     route_ci : in std_logic;
     f0_load : in std_logic;
     f1_load : in std_logic;
     d0_load : in std_logic;
     d1_load : in std_logic;
     ce0 : out std_logic;
     cl0 : out std_logic;
     z0 : out std_logic;
     ff0 : out std_logic;
     ce1 : out std_logic;
     cl1 : out std_logic;
     z1 : out std_logic;
     ff1 : out std_logic;
     ov_msb : out std_logic;
     co_msb : out std_logic;
     cmsb : out std_logic;
     so : out std_logic;
     f0_bus_stat : out std_logic;
     f0_blk_stat : out std_logic;
     f1_bus_stat : out std_logic;
     f1_blk_stat : out std_logic;
     ce0_reg : out std_logic;
     cl0_reg : out std_logic;
     z0_reg : out std_logic;
     ff0_reg : out std_logic;
     ce1_reg : out std_logic;
     cl1_reg : out std_logic;
     z1_reg : out std_logic;
     ff1_reg : out std_logic;
     ov_msb_reg : out std_logic;
     co_msb_reg : out std_logic;
     cmsb_reg : out std_logic;
     so_reg : out std_logic;
     f0_bus_stat_reg : out std_logic;
     f0_blk_stat_reg : out std_logic;
     f1_bus_stat_reg : out std_logic;
     f1_blk_stat_reg : out std_logic);

end component;
component cy_psoc3_dp16
    generic(cy_dpconfig_a : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     cy_dpconfig_b : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_b : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_b : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_b : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_b : std_logic_vector (7 downto 0) := (others => '0');
     ce0_sync : std_logic_vector (1 downto 0) := (others => '1');
     cl0_sync : std_logic_vector (1 downto 0) := (others => '1');
     z0_sync : std_logic_vector (1 downto 0) := (others => '1');
     ff0_sync : std_logic_vector (1 downto 0) := (others => '1');
     ce1_sync : std_logic_vector (1 downto 0) := (others => '1');
     cl1_sync : std_logic_vector (1 downto 0) := (others => '1');
     z1_sync : std_logic_vector (1 downto 0) := (others => '1');
     ff1_sync : std_logic_vector (1 downto 0) := (others => '1');
     ov_msb_sync : std_logic_vector (1 downto 0) := (others => '1');
     co_msb_sync : std_logic_vector (1 downto 0) := (others => '1');
     cmsb_sync : std_logic_vector (1 downto 0) := (others => '1');
     so_sync : std_logic_vector (1 downto 0) := (others => '1');
     f0_bus_sync : std_logic_vector (1 downto 0) := (others => '1');
     f0_blk_sync : std_logic_vector (1 downto 0) := (others => '1');
     f1_bus_sync : std_logic_vector (1 downto 0) := (others => '1');
     f1_blk_sync : std_logic_vector (1 downto 0) := (others => '1'));
    port ( reset : in std_logic := '0';
     clk : in std_logic;
     cs_addr : in std_logic_vector (2 downto 0);
     route_si : in std_logic;
     route_ci : in std_logic;
     f0_load : in std_logic;
     f1_load : in std_logic;
     d0_load : in std_logic;
     d1_load : in std_logic;
     ce0 : out std_logic_vector (1 downto 0);
     cl0 : out std_logic_vector (1 downto 0);
     z0 : out std_logic_vector (1 downto 0);
     ff0 : out std_logic_vector (1 downto 0);
     ce1 : out std_logic_vector (1 downto 0);
     cl1 : out std_logic_vector (1 downto 0);
     z1 : out std_logic_vector (1 downto 0);
     ff1 : out std_logic_vector (1 downto 0);
     ov_msb : out std_logic_vector (1 downto 0);
     co_msb : out std_logic_vector (1 downto 0);
     cmsb : out std_logic_vector (1 downto 0);
     so : out std_logic_vector (1 downto 0);
     f0_bus_stat : out std_logic_vector (1 downto 0);
     f0_blk_stat : out std_logic_vector (1 downto 0);
     f1_bus_stat : out std_logic_vector (1 downto 0);
     f1_blk_stat : out std_logic_vector (1 downto 0);
     ce0_reg : out std_logic_vector (1 downto 0);
     cl0_reg : out std_logic_vector (1 downto 0);
     z0_reg : out std_logic_vector (1 downto 0);
     ff0_reg : out std_logic_vector (1 downto 0);
     ce1_reg : out std_logic_vector (1 downto 0);
     cl1_reg : out std_logic_vector (1 downto 0);
     z1_reg : out std_logic_vector (1 downto 0);
     ff1_reg : out std_logic_vector (1 downto 0);
     ov_msb_reg : out std_logic_vector (1 downto 0);
     co_msb_reg : out std_logic_vector (1 downto 0);
     cmsb_reg : out std_logic_vector (1 downto 0);
     so_reg : out std_logic_vector (1 downto 0);
     f0_bus_stat_reg : out std_logic_vector (1 downto 0);
     f0_blk_stat_reg : out std_logic_vector (1 downto 0);
     f1_bus_stat_reg : out std_logic_vector (1 downto 0);
     f1_blk_stat_reg : out std_logic_vector (1 downto 0));
end component;
component cy_psoc3_dp24
    generic(cy_dpconfig_a : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     cy_dpconfig_b : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_b : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_b : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_b : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_b : std_logic_vector (7 downto 0) := (others => '0');
     cy_dpconfig_c : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_c : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_c : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_c : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_c : std_logic_vector (7 downto 0) := (others => '0');
     ce0_sync : std_logic_vector (2 downto 0) := (others => '1');
     cl0_sync : std_logic_vector (2 downto 0) := (others => '1');
     z0_sync : std_logic_vector (2 downto 0) := (others => '1');
     ff0_sync : std_logic_vector (2 downto 0) := (others => '1');
     ce1_sync : std_logic_vector (2 downto 0) := (others => '1');
     cl1_sync : std_logic_vector (2 downto 0) := (others => '1');
     z1_sync : std_logic_vector (2 downto 0) := (others => '1');
     ff1_sync : std_logic_vector (2 downto 0) := (others => '1');
     ov_msb_sync : std_logic_vector (2 downto 0) := (others => '1');
     co_msb_sync : std_logic_vector (2 downto 0) := (others => '1');
     cmsb_sync : std_logic_vector (2 downto 0) := (others => '1');
     so_sync : std_logic_vector (2 downto 0) := (others => '1');
     f0_bus_sync : std_logic_vector (2 downto 0) := (others => '1');
     f0_blk_sync : std_logic_vector (2 downto 0) := (others => '1');
     f1_bus_sync : std_logic_vector (2 downto 0) := (others => '1');
     f1_blk_sync : std_logic_vector (2 downto 0) := (others => '1'));
    port ( reset : in std_logic := '0';
     clk : in std_logic;
     cs_addr : in std_logic_vector (2 downto 0);
     route_si : in std_logic;
     route_ci : in std_logic;
     f0_load : in std_logic;
     f1_load : in std_logic;
     d0_load : in std_logic;
     d1_load : in std_logic;
     ce0 : out std_logic_vector (2 downto 0);
     cl0 : out std_logic_vector (2 downto 0);
     z0 : out std_logic_vector (2 downto 0);
     ff0 : out std_logic_vector (2 downto 0);
     ce1 : out std_logic_vector (2 downto 0);
     cl1 : out std_logic_vector (2 downto 0);
     z1 : out std_logic_vector (2 downto 0);
     ff1 : out std_logic_vector (2 downto 0);
     ov_msb : out std_logic_vector (2 downto 0);
     co_msb : out std_logic_vector (2 downto 0);
     cmsb : out std_logic_vector (2 downto 0);
     so : out std_logic_vector (2 downto 0);
     f0_bus_stat : out std_logic_vector (2 downto 0);
     f0_blk_stat : out std_logic_vector (2 downto 0);
     f1_bus_stat : out std_logic_vector (2 downto 0);
     f1_blk_stat : out std_logic_vector (2 downto 0);
     ce0_reg : out std_logic_vector (2 downto 0);
     cl0_reg : out std_logic_vector (2 downto 0);
     z0_reg : out std_logic_vector (2 downto 0);
     ff0_reg : out std_logic_vector (2 downto 0);
     ce1_reg : out std_logic_vector (2 downto 0);
     cl1_reg : out std_logic_vector (2 downto 0);
     z1_reg : out std_logic_vector (2 downto 0);
     ff1_reg : out std_logic_vector (2 downto 0);
     ov_msb_reg : out std_logic_vector (2 downto 0);
     co_msb_reg : out std_logic_vector (2 downto 0);
     cmsb_reg : out std_logic_vector (2 downto 0);
     so_reg : out std_logic_vector (2 downto 0);
     f0_bus_stat_reg : out std_logic_vector (2 downto 0);
     f0_blk_stat_reg : out std_logic_vector (2 downto 0);
     f1_bus_stat_reg : out std_logic_vector (2 downto 0);
     f1_blk_stat_reg : out std_logic_vector (2 downto 0));
end component;
component cy_psoc3_dp32
    generic(cy_dpconfig_a : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_a : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_a : std_logic_vector (7 downto 0) := (others => '0');
     cy_dpconfig_b : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_b : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_b : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_b : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_b : std_logic_vector (7 downto 0) := (others => '0');
     cy_dpconfig_c : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_c : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_c : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_c : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_c : std_logic_vector (7 downto 0) := (others => '0');
     cy_dpconfig_d : std_logic_vector (207 downto 0) :=
     X"0000_0000_0000_0000_0000_0000_0000_0000_FFFF_FFFF_0000_0000_0000";
     d0_init_d : std_logic_vector (7 downto 0) := (others => '0');
     d1_init_d : std_logic_vector (7 downto 0) := (others => '0');
     a0_init_d : std_logic_vector (7 downto 0) := (others => '0');
     a1_init_d : std_logic_vector (7 downto 0) := (others => '0');
     ce0_sync : std_logic_vector (3 downto 0) := (others => '1');
     cl0_sync : std_logic_vector (3 downto 0) := (others => '1');
     z0_sync : std_logic_vector (3 downto 0) := (others => '1');
     ff0_sync : std_logic_vector (3 downto 0) := (others => '1');
     ce1_sync : std_logic_vector (3 downto 0) := (others => '1');
     cl1_sync : std_logic_vector (3 downto 0) := (others => '1');
     z1_sync : std_logic_vector (3 downto 0) := (others => '1');
     ff1_sync : std_logic_vector (3 downto 0) := (others => '1');
     ov_msb_sync : std_logic_vector (3 downto 0) := (others => '1');
     co_msb_sync : std_logic_vector (3 downto 0) := (others => '1');
     cmsb_sync : std_logic_vector (3 downto 0) := (others => '1');
     so_sync : std_logic_vector (3 downto 0) := (others => '1');
     f0_bus_sync : std_logic_vector (3 downto 0) := (others => '1');
     f0_blk_sync : std_logic_vector (3 downto 0) := (others => '1');
     f1_bus_sync : std_logic_vector (3 downto 0) := (others => '1');
     f1_blk_sync : std_logic_vector (3 downto 0) := (others => '1'));
    port ( reset : in std_logic := '0';
     clk : in std_logic;
     cs_addr : in std_logic_vector (2 downto 0);
     route_si : in std_logic;
     route_ci : in std_logic;
     f0_load : in std_logic;
     f1_load : in std_logic;
     d0_load : in std_logic;
     d1_load : in std_logic;
     ce0 : out std_logic_vector (3 downto 0);
     cl0 : out std_logic_vector (3 downto 0);
     z0 : out std_logic_vector (3 downto 0);
     ff0 : out std_logic_vector (3 downto 0);
     ce1 : out std_logic_vector (3 downto 0);
     cl1 : out std_logic_vector (3 downto 0);
     z1 : out std_logic_vector (3 downto 0);
     ff1 : out std_logic_vector (3 downto 0);
     ov_msb : out std_logic_vector (3 downto 0);
     co_msb : out std_logic_vector (3 downto 0);
     cmsb : out std_logic_vector (3 downto 0);
     so : out std_logic_vector (3 downto 0);
     f0_bus_stat : out std_logic_vector (3 downto 0);
     f0_blk_stat : out std_logic_vector (3 downto 0);
     f1_bus_stat : out std_logic_vector (3 downto 0);
     f1_blk_stat : out std_logic_vector (3 downto 0);
     ce0_reg : out std_logic_vector (3 downto 0);
     cl0_reg : out std_logic_vector (3 downto 0);
     z0_reg : out std_logic_vector (3 downto 0);
     ff0_reg : out std_logic_vector (3 downto 0);
     ce1_reg : out std_logic_vector (3 downto 0);
     cl1_reg : out std_logic_vector (3 downto 0);
     z1_reg : out std_logic_vector (3 downto 0);
     ff1_reg : out std_logic_vector (3 downto 0);
     ov_msb_reg : out std_logic_vector (3 downto 0);
     co_msb_reg : out std_logic_vector (3 downto 0);
     cmsb_reg : out std_logic_vector (3 downto 0);
     so_reg : out std_logic_vector (3 downto 0);
     f0_bus_stat_reg : out std_logic_vector (3 downto 0);
     f0_blk_stat_reg : out std_logic_vector (3 downto 0);
     f1_bus_stat_reg : out std_logic_vector (3 downto 0);
     f1_blk_stat_reg : out std_logic_vector (3 downto 0));
end component;
component cy_psoc3_control_wrapper
    generic(cy_force_order : boolean := false);
    port (control : out std_logic_vector (7 downto 0));
end component;

end psoc3pkg;

package body psoc3pkg is
end psoc3pkg;
